


module exp_const(output logic y,
                 input logic clk, n_rst);

parameter OFFSET = 0;


// e ^ -2
// logic [1023:0] exp_value = 1023'b00000000010000100001010000000000010000000000010000000000000100001000000000000000000100001000001000000000100000100100000010100000000000000000000000000101000000010100000000000000000100101000001000000001101000000000100000010011100010000001000010000000001000000001000000010000001000011000000100000000000000000000100000110100001000100000000000000000000000000000010001010000001000000000000000000001001000010100100000100000000000000000010010000101001000001000000000000010000000000000000000000000000110010000000000000000001110010000100000000000100000000000100000000000000000000000000000000000000000001000111000000000000010010000001000000000100000110000110010000010010000000000000000000000000000111000001000001000100110000000010010000100000000000000000000000001000000100000001000000000000100100000000000010000100100000000001000100000101000000000000000000000000001000000000000010000000000000000001000000000000100000000000000000000000000000100000000000001000100000001000000100100000000001100010000001000000100100001110000010001000000000001010000000100001000000000000000100001001000000101100000000000010010100000;

// e ^ -4
logic [1023:0] exp_value = 1023'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100010000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000;

int i = 0;

assign y = exp_value[i];

always_ff @(posedge clk, negedge n_rst) begin
    if(~n_rst)
        i <= OFFSET;
    else 
        i <= (i + 1) % 1024;
end

endmodule