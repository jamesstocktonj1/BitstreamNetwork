`timescale 1ns / 1ps


module network_tb;

const int bitstream_length = 256;

logic clk, n_rst, compute;

int x [0:1];
int y [0:0];

int i = 0;
int j = 0;
int k = 0;

int dataFile;


int points_data1 [0:249] = {
	129,
	93,
	55,
	120,
	137,
	149,
	180,
	119,
	104,
	86,
	66,
	79,
	125,
	84,
	155,
	138,
	79,
	141,
	211,
	88,
	133,
	107,
	141,
	84,
	135,
	107,
	96,
	107,
	87,
	201,
	83,
	102,
	60,
	120,
	129,
	98,
	163,
	80,
	163,
	134,
	78,
	161,
	114,
	159,
	70,
	166,
	78,
	97,
	142,
	54,
	140,
	67,
	62,
	97,
	172,
	172,
	84,
	113,
	52,
	74,
	144,
	175,
	0,
	63,
	95,
	104,
	88,
	98,
	129,
	159,
	69,
	93,
	140,
	157,
	85,
	45,
	64,
	203,
	64,
	120,
	153,
	131,
	75,
	145,
	96,
	92,
	75,
	143,
	171,
	89,
	109,
	91,
	60,
	124,
	120,
	151,
	81,
	68,
	164,
	135,
	112,
	164,
	67,
	135,
	131,
	118,
	89,
	124,
	109,
	152,
	130,
	112,
	145,
	86,
	132,
	118,
	85,
	171,
	15,
	152,
	133,
	112,
	94,
	151,
	117,
	185,
	220,
	179,
	206,
	204,
	209,
	162,
	185,
	122,
	203,
	176,
	170,
	192,
	137,
	238,
	129,
	105,
	193,
	120,
	240,
	197,
	173,
	182,
	175,
	162,
	148,
	175,
	230,
	164,
	141,
	122,
	184,
	184,
	166,
	158,
	165,
	241,
	174,
	214,
	211,
	193,
	224,
	183,
	198,
	224,
	205,
	186,
	178,
	169,
	78,
	137,
	193,
	256,
	197,
	160,
	198,
	215,
	230,
	185,
	150,
	100,
	147,
	202,
	168,
	115,
	108,
	175,
	130,
	190,
	206,
	233,
	139,
	238,
	146,
	231,
	160,
	207,
	149,
	96,
	161,
	227,
	181,
	203,
	215,
	251,
	173,
	152,
	231,
	197,
	128,
	187,
	151,
	115,
	150,
	110,
	218,
	151,
	161,
	136,
	176,
	191,
	198,
	178,
	156,
	144,
	181,
	141,
	170,
	177,
	214,
	208,
	196,
	168,
	198,
	202,
	185,
	179,
	175,
	189,
	165,
	78,
	161,
	187,
	185,
	94
};

int points_data2 [0:249] = {
	105,
	151,
	141,
	102,
	103,
	107,
	100,
	100,
	126,
	155,
	126,
	155,
	77,
	110,
	79,
	125,
	116,
	120,
	56,
	127,
	110,
	114,
	88,
	149,
	86,
	120,
	148,
	110,
	119,
	91,
	114,
	115,
	138,
	120,
	110,
	113,
	132,
	117,
	106,
	95,
	107,
	106,
	96,
	109,
	116,
	86,
	117,
	143,
	121,
	127,
	117,
	132,
	124,
	108,
	96,
	81,
	123,
	108,
	113,
	118,
	122,
	103,
	165,
	131,
	103,
	112,
	116,
	123,
	93,
	107,
	123,
	133,
	81,
	101,
	145,
	127,
	100,
	115,
	120,
	144,
	137,
	98,
	110,
	118,
	110,
	129,
	130,
	89,
	103,
	149,
	98,
	104,
	130,
	125,
	117,
	101,
	111,
	119,
	121,
	123,
	106,
	109,
	120,
	102,
	68,
	119,
	123,
	122,
	112,
	114,
	118,
	146,
	129,
	111,
	117,
	128,
	153,
	104,
	132,
	138,
	107,
	100,
	139,
	112,
	129,
	192,
	165,
	181,
	184,
	166,
	153,
	188,
	155,
	193,
	163,
	158,
	185,
	210,
	202,
	185,
	201,
	216,
	166,
	186,
	158,
	190,
	179,
	193,
	180,
	164,
	188,
	194,
	179,
	179,
	185,
	181,
	154,
	182,
	181,
	185,
	160,
	151,
	194,
	189,
	159,
	170,
	167,
	165,
	174,
	178,
	157,
	172,
	179,
	179,
	248,
	179,
	163,
	167,
	163,
	167,
	186,
	166,
	180,
	192,
	152,
	199,
	196,
	182,
	163,
	211,
	196,
	158,
	192,
	186,
	161,
	175,
	182,
	168,
	167,
	123,
	166,
	150,
	180,
	214,
	209,
	150,
	156,
	190,
	170,
	162,
	174,
	163,
	164,
	170,
	204,
	162,
	198,
	177,
	182,
	194,
	203,
	172,
	175,
	188,
	176,
	163,
	150,
	194,
	205,
	172,
	160,
	211,
	161,
	175,
	176,
	164,
	141,
	178,
	206,
	198,
	187,
	175,
	181,
	184,
	160,
	219,
	199,
	171,
	178,
	215
};

int data_perceptron1 [0:249] = {
	107,
	103,
	95,
	138,
	120,
	107,
	12,
	101,
	164,
	139,
	171,
	154,
	159,
	58,
	40,
	131,
	140,
	97,
	107,
	125,
	109,
	122,
	48,
	126,
	103,
	110,
	111,
	90,
	161,
	107,
	95,
	120,
	0,
	103,
	214,
	48,
	62,
	135,
	94,
	177,
	125,
	145,
	75,
	57,
	136,
	103,
	113,
	27,
	90,
	170,
	176,
	90,
	98,
	142,
	84,
	151,
	53,
	112,
	38,
	159,
	141,
	79,
	50,
	122,
	77,
	58,
	136,
	66,
	64,
	149,
	124,
	105,
	116,
	103,
	204,
	65,
	110,
	147,
	93,
	178,
	99,
	95,
	81,
	152,
	78,
	105,
	45,
	131,
	162,
	154,
	103,
	105,
	96,
	81,
	93,
	142,
	125,
	135,
	59,
	90,
	57,
	158,
	67,
	181,
	111,
	38,
	102,
	90,
	86,
	94,
	157,
	99,
	125,
	87,
	88,
	135,
	143,
	76,
	81,
	81,
	74,
	97,
	23,
	135,
	113,
	171,
	156,
	123,
	190,
	182,
	165,
	145,
	183,
	144,
	198,
	214,
	145,
	212,
	214,
	62,
	217,
	202,
	105,
	211,
	181,
	170,
	215,
	218,
	147,
	185,
	179,
	148,
	226,
	181,
	157,
	90,
	200,
	222,
	171,
	254,
	151,
	153,
	153,
	173,
	53,
	97,
	118,
	172,
	107,
	149,
	154,
	176,
	179,
	199,
	232,
	179,
	176,
	90,
	225,
	226,
	196,
	182,
	163,
	140,
	216,
	147,
	134,
	184,
	204,
	191,
	186,
	173,
	123,
	139,
	159,
	120,
	141,
	177,
	152,
	160,
	138,
	173,
	178,
	209,
	158,
	185,
	111,
	120,
	236,
	191,
	144,
	80,
	96,
	185,
	160,
	143,
	153,
	161,
	100,
	153,
	179,
	178,
	141,
	190,
	169,
	199,
	103,
	180,
	99,
	188,
	176,
	192,
	180,
	137,
	180,
	172,
	129,
	256,
	170,
	140,
	193,
	140,
	149,
	154,
	96,
	96,
	153,
	186,
	132,
	132
};

int data_perceptron2 [0:249] = {
	89,
	83,
	104,
	115,
	85,
	105,
	159,
	93,
	101,
	115,
	85,
	94,
	67,
	113,
	126,
	77,
	87,
	91,
	112,
	81,
	96,
	97,
	134,
	114,
	125,
	107,
	100,
	91,
	84,
	94,
	120,
	74,
	145,
	93,
	79,
	144,
	155,
	108,
	120,
	60,
	109,
	95,
	93,
	105,
	87,
	103,
	104,
	120,
	107,
	100,
	51,
	109,
	125,
	79,
	106,
	64,
	112,
	73,
	147,
	100,
	94,
	120,
	114,
	84,
	104,
	112,
	95,
	125,
	108,
	93,
	106,
	108,
	109,
	101,
	48,
	100,
	93,
	92,
	110,
	97,
	109,
	92,
	117,
	108,
	117,
	97,
	119,
	82,
	74,
	84,
	92,
	101,
	90,
	112,
	106,
	102,
	90,
	127,
	119,
	101,
	109,
	102,
	89,
	71,
	99,
	134,
	99,
	113,
	103,
	124,
	74,
	129,
	84,
	136,
	114,
	81,
	75,
	128,
	124,
	128,
	108,
	113,
	121,
	84,
	129,
	149,
	154,
	159,
	133,
	154,
	166,
	159,
	193,
	157,
	175,
	179,
	156,
	148,
	142,
	205,
	146,
	151,
	206,
	155,
	163,
	157,
	166,
	146,
	159,
	152,
	147,
	164,
	152,
	151,
	171,
	174,
	179,
	147,
	164,
	129,
	158,
	153,
	181,
	168,
	193,
	202,
	182,
	147,
	169,
	177,
	157,
	149,
	119,
	153,
	119,
	163,
	185,
	196,
	146,
	139,
	167,
	156,
	166,
	195,
	147,
	128,
	164,
	142,
	135,
	170,
	147,
	157,
	189,
	159,
	149,
	169,
	169,
	141,
	155,
	156,
	161,
	169,
	171,
	165,
	181,
	163,
	175,
	188,
	151,
	152,
	175,
	189,
	176,
	141,
	140,
	141,
	168,
	144,
	183,
	198,
	162,
	169,
	164,
	166,
	160,
	138,
	181,
	150,
	168,
	163,
	175,
	182,
	152,
	179,
	142,
	182,
	193,
	122,
	147,
	147,
	168,
	171,
	185,
	174,
	203,
	182,
	191,
	137,
	202,
	170
};


// assign x[0] = j * 5;
// assign x[1] = k * 5;

assign x[0] = data_perceptron1[j];
assign x[1] = data_perceptron2[j];

network n(
    .clk(clk),
    .n_rst(n_rst),
	.compute(compute),
    .network_input(x),
    .network_output(y)
);
defparam n.SEED = 8'b10001101;


initial begin
    dataFile = $fopen("data/log.txt", "w");

    clk = 1'b0;
    n_rst = 1'b1;
	compute = 1'b0;

    #20ps n_rst = 1'b0;
    #20ps n_rst = 1'b1;


	for(j=0; j<250; j++) begin
		compute = 1'b1;

		for(i=0; i<bitstream_length; i++) begin
			#10ps clk = ~clk;
			#10ps clk = ~clk;
		end

		compute = 1'b0;
		#10ps clk = ~clk;
		#10ps clk = ~clk;

			$fwrite(dataFile, "%f\n", real'(y[0])/bitstream_length);
	end

    $fclose();
    $stop();
end

endmodule