`timescale 1ns / 1ps


module network_tb;

logic x1;
logic x2;
logic [1:0] x;
logic y;
logic clk;
logic n_rst;

int i = 0;
int j = 0;
int k = 0;

real val = 0.0;
real value = 0.0;

int dataFile;


int points_data1 [0:249] = {
	129,
	93,
	55,
	120,
	137,
	149,
	180,
	119,
	104,
	86,
	66,
	79,
	125,
	84,
	155,
	138,
	79,
	141,
	211,
	88,
	133,
	107,
	141,
	84,
	135,
	107,
	96,
	107,
	87,
	201,
	83,
	102,
	60,
	120,
	129,
	98,
	163,
	80,
	163,
	134,
	78,
	161,
	114,
	159,
	70,
	166,
	78,
	97,
	142,
	54,
	140,
	67,
	62,
	97,
	172,
	172,
	84,
	113,
	52,
	74,
	144,
	175,
	0,
	63,
	95,
	104,
	88,
	98,
	129,
	159,
	69,
	93,
	140,
	157,
	85,
	45,
	64,
	203,
	64,
	120,
	153,
	131,
	75,
	145,
	96,
	92,
	75,
	143,
	171,
	89,
	109,
	91,
	60,
	124,
	120,
	151,
	81,
	68,
	164,
	135,
	112,
	164,
	67,
	135,
	131,
	118,
	89,
	124,
	109,
	152,
	130,
	112,
	145,
	86,
	132,
	118,
	85,
	171,
	15,
	152,
	133,
	112,
	94,
	151,
	117,
	185,
	220,
	179,
	206,
	204,
	209,
	162,
	185,
	122,
	203,
	176,
	170,
	192,
	137,
	238,
	129,
	105,
	193,
	120,
	240,
	197,
	173,
	182,
	175,
	162,
	148,
	175,
	230,
	164,
	141,
	122,
	184,
	184,
	166,
	158,
	165,
	241,
	174,
	214,
	211,
	193,
	224,
	183,
	198,
	224,
	205,
	186,
	178,
	169,
	78,
	137,
	193,
	256,
	197,
	160,
	198,
	215,
	230,
	185,
	150,
	100,
	147,
	202,
	168,
	115,
	108,
	175,
	130,
	190,
	206,
	233,
	139,
	238,
	146,
	231,
	160,
	207,
	149,
	96,
	161,
	227,
	181,
	203,
	215,
	251,
	173,
	152,
	231,
	197,
	128,
	187,
	151,
	115,
	150,
	110,
	218,
	151,
	161,
	136,
	176,
	191,
	198,
	178,
	156,
	144,
	181,
	141,
	170,
	177,
	214,
	208,
	196,
	168,
	198,
	202,
	185,
	179,
	175,
	189,
	165,
	78,
	161,
	187,
	185,
	94
};

int points_data2 [0:249] = {
	105,
	151,
	141,
	102,
	103,
	107,
	100,
	100,
	126,
	155,
	126,
	155,
	77,
	110,
	79,
	125,
	116,
	120,
	56,
	127,
	110,
	114,
	88,
	149,
	86,
	120,
	148,
	110,
	119,
	91,
	114,
	115,
	138,
	120,
	110,
	113,
	132,
	117,
	106,
	95,
	107,
	106,
	96,
	109,
	116,
	86,
	117,
	143,
	121,
	127,
	117,
	132,
	124,
	108,
	96,
	81,
	123,
	108,
	113,
	118,
	122,
	103,
	165,
	131,
	103,
	112,
	116,
	123,
	93,
	107,
	123,
	133,
	81,
	101,
	145,
	127,
	100,
	115,
	120,
	144,
	137,
	98,
	110,
	118,
	110,
	129,
	130,
	89,
	103,
	149,
	98,
	104,
	130,
	125,
	117,
	101,
	111,
	119,
	121,
	123,
	106,
	109,
	120,
	102,
	68,
	119,
	123,
	122,
	112,
	114,
	118,
	146,
	129,
	111,
	117,
	128,
	153,
	104,
	132,
	138,
	107,
	100,
	139,
	112,
	129,
	192,
	165,
	181,
	184,
	166,
	153,
	188,
	155,
	193,
	163,
	158,
	185,
	210,
	202,
	185,
	201,
	216,
	166,
	186,
	158,
	190,
	179,
	193,
	180,
	164,
	188,
	194,
	179,
	179,
	185,
	181,
	154,
	182,
	181,
	185,
	160,
	151,
	194,
	189,
	159,
	170,
	167,
	165,
	174,
	178,
	157,
	172,
	179,
	179,
	248,
	179,
	163,
	167,
	163,
	167,
	186,
	166,
	180,
	192,
	152,
	199,
	196,
	182,
	163,
	211,
	196,
	158,
	192,
	186,
	161,
	175,
	182,
	168,
	167,
	123,
	166,
	150,
	180,
	214,
	209,
	150,
	156,
	190,
	170,
	162,
	174,
	163,
	164,
	170,
	204,
	162,
	198,
	177,
	182,
	194,
	203,
	172,
	175,
	188,
	176,
	163,
	150,
	194,
	205,
	172,
	160,
	211,
	161,
	175,
	176,
	164,
	141,
	178,
	206,
	198,
	187,
	175,
	181,
	184,
	160,
	219,
	199,
	171,
	178,
	215
};


generator x1_gen(
	.clk(clk),
	.n_rst(n_rst),
	.x(j * 5),
	.y(x1)
);
// defparam x1_gen.SEED = 0'b101010;

generator x2_gen(
	.clk(clk),
	.n_rst(n_rst),
	.x(k * 5),
	.y(x2)
);

assign x = {x1, x2};

network n(
    .clk(clk),
    .n_rst(n_rst),
    .network_input(x),
    .network_output(y)
);


initial begin
    dataFile = $fopen("data/log.txt", "w");

    clk = 1'b0;
    n_rst = 1'b1;

    #20ps n_rst = 1'b0;
    #20ps n_rst = 1'b1;
end

always #10ps clk = ~clk;


always_ff @(posedge clk) begin

    if(i < 256) begin
        i++;
        if(y)
            value++;
    end
    else begin
        val <= real'(value / 256);
        $fwrite(dataFile, "%f\n", val);

        i <= 0;
        value <= 0.0;

        if(j < 49)
            j++;
        else begin
			j <= 0;
			if(k < 49)
				k++;
			else begin
				$fclose(dataFile);
            	$stop();
			end
        end
    end
end

endmodule