`timescale 1ns / 1ps


module network_tb;

const int bitstream_length = 256;

logic clk, n_rst, compute;

int x [0:1];
int y [0:0];

int i = 0;
int j = 0;
int k = 0;

int dataFile;


int data_perceptron1 [0:249] = {
	107,
	103,
	95,
	138,
	120,
	107,
	12,
	101,
	164,
	139,
	171,
	154,
	159,
	58,
	40,
	131,
	140,
	97,
	107,
	125,
	109,
	122,
	48,
	126,
	103,
	110,
	111,
	90,
	161,
	107,
	95,
	120,
	0,
	103,
	214,
	48,
	62,
	135,
	94,
	177,
	125,
	145,
	75,
	57,
	136,
	103,
	113,
	27,
	90,
	170,
	176,
	90,
	98,
	142,
	84,
	151,
	53,
	112,
	38,
	159,
	141,
	79,
	50,
	122,
	77,
	58,
	136,
	66,
	64,
	149,
	124,
	105,
	116,
	103,
	204,
	65,
	110,
	147,
	93,
	178,
	99,
	95,
	81,
	152,
	78,
	105,
	45,
	131,
	162,
	154,
	103,
	105,
	96,
	81,
	93,
	142,
	125,
	135,
	59,
	90,
	57,
	158,
	67,
	181,
	111,
	38,
	102,
	90,
	86,
	94,
	157,
	99,
	125,
	87,
	88,
	135,
	143,
	76,
	81,
	81,
	74,
	97,
	23,
	135,
	113,
	171,
	156,
	123,
	190,
	182,
	165,
	145,
	183,
	144,
	198,
	214,
	145,
	212,
	214,
	62,
	217,
	202,
	105,
	211,
	181,
	170,
	215,
	218,
	147,
	185,
	179,
	148,
	226,
	181,
	157,
	90,
	200,
	222,
	171,
	254,
	151,
	153,
	153,
	173,
	53,
	97,
	118,
	172,
	107,
	149,
	154,
	176,
	179,
	199,
	232,
	179,
	176,
	90,
	225,
	226,
	196,
	182,
	163,
	140,
	216,
	147,
	134,
	184,
	204,
	191,
	186,
	173,
	123,
	139,
	159,
	120,
	141,
	177,
	152,
	160,
	138,
	173,
	178,
	209,
	158,
	185,
	111,
	120,
	236,
	191,
	144,
	80,
	96,
	185,
	160,
	143,
	153,
	161,
	100,
	153,
	179,
	178,
	141,
	190,
	169,
	199,
	103,
	180,
	99,
	188,
	176,
	192,
	180,
	137,
	180,
	172,
	129,
	256,
	170,
	140,
	193,
	140,
	149,
	154,
	96,
	96,
	153,
	186,
	132,
	132
};

int data_perceptron2 [0:249] = {
	89,
	83,
	104,
	115,
	85,
	105,
	159,
	93,
	101,
	115,
	85,
	94,
	67,
	113,
	126,
	77,
	87,
	91,
	112,
	81,
	96,
	97,
	134,
	114,
	125,
	107,
	100,
	91,
	84,
	94,
	120,
	74,
	145,
	93,
	79,
	144,
	155,
	108,
	120,
	60,
	109,
	95,
	93,
	105,
	87,
	103,
	104,
	120,
	107,
	100,
	51,
	109,
	125,
	79,
	106,
	64,
	112,
	73,
	147,
	100,
	94,
	120,
	114,
	84,
	104,
	112,
	95,
	125,
	108,
	93,
	106,
	108,
	109,
	101,
	48,
	100,
	93,
	92,
	110,
	97,
	109,
	92,
	117,
	108,
	117,
	97,
	119,
	82,
	74,
	84,
	92,
	101,
	90,
	112,
	106,
	102,
	90,
	127,
	119,
	101,
	109,
	102,
	89,
	71,
	99,
	134,
	99,
	113,
	103,
	124,
	74,
	129,
	84,
	136,
	114,
	81,
	75,
	128,
	124,
	128,
	108,
	113,
	121,
	84,
	129,
	149,
	154,
	159,
	133,
	154,
	166,
	159,
	193,
	157,
	175,
	179,
	156,
	148,
	142,
	205,
	146,
	151,
	206,
	155,
	163,
	157,
	166,
	146,
	159,
	152,
	147,
	164,
	152,
	151,
	171,
	174,
	179,
	147,
	164,
	129,
	158,
	153,
	181,
	168,
	193,
	202,
	182,
	147,
	169,
	177,
	157,
	149,
	119,
	153,
	119,
	163,
	185,
	196,
	146,
	139,
	167,
	156,
	166,
	195,
	147,
	128,
	164,
	142,
	135,
	170,
	147,
	157,
	189,
	159,
	149,
	169,
	169,
	141,
	155,
	156,
	161,
	169,
	171,
	165,
	181,
	163,
	175,
	188,
	151,
	152,
	175,
	189,
	176,
	141,
	140,
	141,
	168,
	144,
	183,
	198,
	162,
	169,
	164,
	166,
	160,
	138,
	181,
	150,
	168,
	163,
	175,
	182,
	152,
	179,
	142,
	182,
	193,
	122,
	147,
	147,
	168,
	171,
	185,
	174,
	203,
	182,
	191,
	137,
	202,
	170
};

int iris_data [0:149][0:3] = {
	{165, 204,  52,  20},
	{159, 175,  52,  20},
	{152, 186,  48,  20},
	{149, 180,  56,  20},
	{162, 209,  52,  20},
	{175, 227,  63,  41},
	{149, 198,  52,  31},
	{162, 198,  56,  20},
	{143, 169,  52,  20},
	{159, 180,  56,  10},
	{175, 215,  56,  20},
	{156, 198,  59,  20},
	{156, 175,  52,  10},
	{139, 175,  41,  10},
	{188, 233,  45,  20},
	{185, 256,  56,  41},
	{175, 227,  48,  41},
	{165, 204,  52,  31},
	{185, 221,  63,  31},
	{165, 221,  56,  31},
	{175, 198,  63,  20},
	{165, 215,  56,  41},
	{149, 209,  37,  20},
	{165, 192,  63,  51},
	{156, 198,  70,  20},
	{162, 175,  59,  20},
	{162, 198,  59,  41},
	{169, 204,  56,  20},
	{169, 198,  52,  20},
	{152, 186,  59,  20},
	{156, 180,  59,  20},
	{175, 198,  56,  41},
	{169, 239,  56,  10},
	{178, 244,  52,  20},
	{159, 180,  56,  20},
	{162, 186,  45,  20},
	{178, 204,  48,  20},
	{159, 209,  52,  10},
	{143, 175,  48,  20},
	{165, 198,  56,  20},
	{162, 204,  48,  31},
	{146, 134,  48,  31},
	{143, 186,  48,  20},
	{162, 204,  59,  61},
	{165, 221,  70,  41},
	{156, 175,  52,  31},
	{165, 221,  59,  20},
	{149, 186,  52,  20},
	{172, 215,  56,  20},
	{162, 192,  52,  20},
	{227, 186, 174, 143},
	{207, 186, 167, 154},
	{224, 180, 182, 154},
	{178, 134, 148, 133},
	{211, 163, 171, 154},
	{185, 163, 167, 133},
	{204, 192, 174, 164},
	{159, 140, 122, 102},
	{214, 169, 171, 133},
	{169, 157, 145, 143},
	{162, 116, 130, 102},
	{191, 175, 156, 154},
	{194, 128, 148, 102},
	{198, 169, 174, 143},
	{181, 169, 134, 133},
	{217, 180, 163, 143},
	{181, 175, 167, 154},
	{188, 157, 152, 102},
	{201, 128, 167, 154},
	{181, 145, 145, 113},
	{191, 186, 178, 184},
	{198, 163, 148, 133},
	{204, 145, 182, 154},
	{198, 163, 174, 123},
	{207, 169, 160, 133},
	{214, 175, 163, 143},
	{220, 163, 178, 143},
	{217, 175, 186, 174},
	{194, 169, 167, 154},
	{185, 151, 130, 102},
	{178, 140, 141, 113},
	{178, 140, 137, 102},
	{188, 157, 145, 123},
	{194, 157, 189, 164},
	{175, 175, 167, 154},
	{194, 198, 167, 164},
	{217, 180, 174, 154},
	{204, 134, 163, 133},
	{181, 175, 152, 133},
	{178, 145, 148, 133},
	{178, 151, 163, 123},
	{198, 175, 171, 143},
	{188, 151, 148, 123},
	{162, 134, 122, 102},
	{181, 157, 156, 133},
	{185, 175, 156, 123},
	{185, 169, 156, 133},
	{201, 169, 160, 133},
	{165, 145, 111, 113},
	{185, 163, 152, 133},
	{204, 192, 223, 256},
	{188, 157, 189, 195},
	{230, 175, 219, 215},
	{204, 169, 208, 184},
	{211, 175, 215, 225},
	{246, 175, 245, 215},
	{159, 145, 167, 174},
	{237, 169, 234, 184},
	{217, 145, 215, 184},
	{233, 209, 226, 256},
	{211, 186, 189, 205},
	{207, 157, 197, 195},
	{220, 175, 204, 215},
	{185, 145, 186, 205},
	{188, 163, 189, 246},
	{207, 186, 197, 236},
	{211, 175, 204, 184},
	{250, 221, 249, 225},
	{250, 151, 256, 236},
	{194, 128, 186, 154},
	{224, 186, 211, 236},
	{181, 163, 182, 205},
	{250, 163, 249, 205},
	{204, 157, 182, 184},
	{217, 192, 211, 215},
	{233, 186, 223, 184},
	{201, 163, 178, 184},
	{198, 175, 182, 184},
	{207, 163, 208, 215},
	{233, 175, 215, 164},
	{240, 163, 226, 195},
	{256, 221, 237, 205},
	{207, 163, 208, 225},
	{204, 163, 189, 154},
	{198, 151, 208, 143},
	{250, 175, 226, 236},
	{204, 198, 208, 246},
	{207, 180, 204, 184},
	{194, 175, 178, 184},
	{224, 180, 200, 215},
	{217, 180, 208, 246},
	{224, 180, 189, 236},
	{188, 157, 189, 195},
	{220, 186, 219, 236},
	{217, 192, 211, 256},
	{217, 175, 193, 236},
	{204, 145, 186, 195},
	{211, 175, 193, 205},
	{201, 198, 200, 236},
	{191, 175, 189, 184}
};


assign x[0] = data_perceptron1[j];
assign x[1] = data_perceptron2[j];

network n(
    .clk(clk),
    .n_rst(n_rst),
	.compute(compute),
    .network_input(x),
    .network_output(y)
);
// defparam n.SEED = 8'b10001101;


initial begin
    dataFile = $fopen("data/separation.txt", "w");

    clk = 1'b0;
    n_rst = 1'b1;
	compute = 1'b0;

    #20ps n_rst = 1'b0;
    #20ps n_rst = 1'b1;


	for(j=0; j<250; j++) begin
		compute = 1'b1;

		for(i=0; i<bitstream_length; i++) begin
			#10ps clk = ~clk;
			#10ps clk = ~clk;
		end

		compute = 1'b0;
		#10ps clk = ~clk;
		#10ps clk = ~clk;

		$fwrite(dataFile, "%f\n", real'(y[0])/bitstream_length);
	end

    $fclose();
    $stop();
end

endmodule