


module constant(output logic a2, a3, a4, a5,
                input logic clk, n_rst);

parameter OFFSET = 0;


int i = 0;

logic [511:0] buffer_a2 = 511'b11011000010000100000111100101101001010101101011010000001000011001011000110100100101011011111001111100100010000110000010101101110111011010101110100111001100001001000110010001111010011011110001011001110101001001011110010011000111000011101101110111011101000011010001001110000000000011010101010010001101011011001000001101011100011110010111101010101011000011100100011110111010111110010110100010000000011111010101100110001110011101001011101010110011011001100101000101111001101111001010100110111100011111101010100000111;
logic [511:0] buffer_a3 = 511'b00001011100000100000000001100000000110010001110001001100000100000000101000000111101110010010100000100000010010110110111100111100010010001100100000011001010000000001101100011000001000100100010010001010110001101010001010101001101000000111100100010101001101001000001010010111100000010001011000000100110000000010000010010001011101100001001100010011111000001010000000010100000010010101001001000000000000111010100001000101000000010100110011000000011100000000010111100001000100100000100100100001010111010111000010000000;
logic [511:0] buffer_a4 = 511'b00000000010001000000010000010010110100000010000000101100010000111000000110100000000000000010100001101000010000001001000001000001000001000000000001011001000000000110001000001010100010000001000010001111000010000101001010011000010000000000010000100100000000010000000000001011001111100111010000011000001100000010111010001010100010000000000100000000000000000000101111000001000000100011001000010001000111000100001010000010000110000000000010000000011000100000000111000001001000100000011111110000010000010000000000101010;
logic [511:0] buffer_a5 = 511'b10001000100000110000001011000010100000001000010000100000001000010100100000000110000000100000100001000000100000000000001000000001101001000000011000100000001000001100001100010000011100100100100010000000000000000000000010000100001001010000000000000000000100100000000000001000000000000000101010110000001001001100000000011100000001000000001010100001000010011100000001000100001010000000010100000000001010000000001100100011001001010000000000000000001011000100000000100001000110000001000100000000000000100010000000000001;

assign a2 = buffer_a2[i];
assign a3 = buffer_a3[i];
assign a4 = buffer_a4[i];
assign a5 = buffer_a5[i];

always_ff @(posedge clk, negedge n_rst) begin
    if (~n_rst)
        i <= OFFSET;
    else
        i <= (i + 1) % 512;
end

endmodule